magic
tech sky130A
magscale 1 2
timestamp 1662126094
<< error_p >>
rect 301 187 497 341
rect 301 182 463 187
rect 497 182 631 187
rect 301 173 309 182
rect 469 154 477 173
<< nwell >>
rect 463 182 497 187
rect 309 173 497 182
rect 309 154 469 173
<< pwell >>
rect -211 -310 211 310
<< nmos >>
rect -15 -100 15 100
<< ndiff >>
rect -73 88 -15 100
rect -73 -88 -61 88
rect -27 -88 -15 88
rect -73 -100 -15 -88
rect 15 88 73 100
rect 15 -88 27 88
rect 61 -88 73 88
rect 15 -100 73 -88
<< ndiffc >>
rect -61 -88 -27 88
rect 27 -88 61 88
<< psubdiff >>
rect -175 240 -79 274
rect 79 240 175 274
rect -175 178 -141 240
rect 141 178 175 240
rect -175 -240 -141 -178
rect 141 -240 175 -178
rect -175 -274 -79 -240
rect 79 -274 175 -240
<< psubdiffcont >>
rect -79 240 79 274
rect -175 -178 -141 178
rect 141 -178 175 178
rect -79 -274 79 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -15 100 15 122
rect -15 -127 15 -100
<< polycont >>
rect -17 138 17 172
<< locali >>
rect -175 240 -79 274
rect 79 240 175 274
rect -175 178 -141 240
rect 141 178 175 240
rect -33 138 -17 172
rect 17 138 33 172
rect -175 -240 -141 -178
rect -61 88 -27 104
rect -61 -240 -27 -88
rect 27 88 61 104
rect 27 -104 61 -88
rect 141 -240 175 -178
rect -175 -274 -79 -240
rect 79 -274 175 -240
rect -823 -908 -622 -856
rect -823 -1008 -763 -908
rect -657 -966 -622 -908
rect -61 -966 -27 -274
rect -657 -1000 -27 -966
rect -657 -1008 -622 -1000
rect -823 -1058 -622 -1008
<< viali >>
rect -17 138 17 172
rect -61 -88 -27 88
rect 27 -88 61 88
rect -763 -1008 -657 -908
<< metal1 >>
rect -7819 3585 -3812 3771
rect -7810 2479 -7641 3585
rect -3998 3167 -3812 3585
rect -3998 2981 -3809 3167
rect -7430 2528 -7290 2544
rect -4000 2528 -3811 2595
rect -7430 2420 -3811 2528
rect -7430 2158 -7290 2420
rect -4000 2393 -3811 2420
rect -7788 2018 -7290 2158
rect -4005 2019 -3816 2039
rect -7105 1863 -3816 2019
rect -7105 1766 -6949 1863
rect -4005 1837 -3816 1863
rect -7796 1610 -6949 1766
rect -4123 1374 -3809 1461
rect -7786 1355 -6164 1356
rect -4124 1355 -3809 1374
rect -7786 1272 -3809 1355
rect -7786 1220 -4170 1272
rect -3998 1259 -3809 1272
rect -7720 844 -6872 878
rect -6906 774 -6872 844
rect -3999 774 -3810 864
rect -6906 740 -1062 774
rect -3999 662 -3810 740
rect -7777 429 -4525 548
rect -4644 276 -4525 429
rect -4001 276 -3812 301
rect -7818 -12 -5017 188
rect -4644 157 -3812 276
rect -4001 99 -3812 157
rect -1096 172 -1062 740
rect -29 172 29 178
rect 289 173 497 187
rect 289 172 469 173
rect -1096 138 -17 172
rect 17 154 469 172
rect 17 138 315 154
rect -29 132 29 138
rect -67 88 -21 100
rect -7818 -412 -5488 -212
rect -5182 -271 -5051 -12
rect -67 -88 -61 88
rect -27 -88 -21 88
rect -67 -100 -21 -88
rect 21 88 67 100
rect 21 -88 27 88
rect 61 -88 67 88
rect 21 -100 67 -88
rect -5182 -290 -3843 -271
rect -5182 -402 -3810 -290
rect 26 -360 60 -100
rect 26 -394 492 -360
rect -7793 -787 -5933 -636
rect -7796 -1190 -6380 -1033
rect -6537 -2476 -6380 -1190
rect -6084 -1449 -5933 -787
rect -5688 -855 -5488 -412
rect -3999 -492 -3810 -402
rect -5690 -899 -5488 -855
rect -5690 -925 -5487 -899
rect -4003 -925 -3809 -857
rect -5690 -945 -3809 -925
rect -823 -908 -622 -856
rect -5690 -1071 -3810 -945
rect -823 -1008 -763 -908
rect -657 -1008 -622 -908
rect -823 -1058 -622 -1008
rect -5690 -1079 -3841 -1071
rect -5690 -1080 -5491 -1079
rect -6084 -1600 -3792 -1449
rect -4002 -1669 -3808 -1600
rect -4001 -2476 -3812 -2036
rect -6537 -2613 -3812 -2476
rect -6537 -2633 -3815 -2613
<< properties >>
string FIXED_BBOX -158 -257 158 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
