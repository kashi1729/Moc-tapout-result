magic
tech sky130A
magscale 1 2
timestamp 1662126094
<< poly >>
rect -1006 866 -806 882
rect -1006 832 -990 866
rect -822 832 -806 866
rect -1006 809 -806 832
rect -1006 456 -806 479
rect -1006 422 -990 456
rect -822 422 -806 456
rect -1006 406 -806 422
rect -1006 286 -806 302
rect -1006 252 -990 286
rect -822 252 -806 286
rect -1006 229 -806 252
rect -1006 -124 -806 -101
rect -1006 -158 -990 -124
rect -822 -158 -806 -124
rect -1006 -174 -806 -158
rect -1006 -294 -806 -278
rect -1006 -328 -990 -294
rect -822 -328 -806 -294
rect -1006 -351 -806 -328
rect -1006 -704 -806 -681
rect -1006 -738 -990 -704
rect -822 -738 -806 -704
rect -1006 -754 -806 -738
rect -1006 -874 -806 -858
rect -1006 -908 -990 -874
rect -822 -908 -806 -874
rect -1006 -931 -806 -908
rect -1006 -1284 -806 -1261
rect -1006 -1318 -990 -1284
rect -822 -1318 -806 -1284
rect -1006 -1334 -806 -1318
rect -1006 -1454 -806 -1438
rect -1006 -1488 -990 -1454
rect -822 -1488 -806 -1454
rect -1006 -1511 -806 -1488
rect -1006 -1864 -806 -1841
rect -1006 -1898 -990 -1864
rect -822 -1898 -806 -1864
rect -1006 -1914 -806 -1898
rect -1006 -2034 -806 -2018
rect -1006 -2068 -990 -2034
rect -822 -2068 -806 -2034
rect -1006 -2091 -806 -2068
rect -1006 -2444 -806 -2421
rect -1006 -2478 -990 -2444
rect -822 -2478 -806 -2444
rect -1006 -2494 -806 -2478
rect -1006 -2614 -806 -2598
rect -1006 -2648 -990 -2614
rect -822 -2648 -806 -2614
rect -1006 -2671 -806 -2648
rect -1006 -3024 -806 -3001
rect -1006 -3058 -990 -3024
rect -822 -3058 -806 -3024
rect -1006 -3074 -806 -3058
rect -1006 -3194 -806 -3178
rect -1006 -3228 -990 -3194
rect -822 -3228 -806 -3194
rect -1006 -3251 -806 -3228
rect -1006 -3604 -806 -3581
rect -1006 -3638 -990 -3604
rect -822 -3638 -806 -3604
rect -1006 -3654 -806 -3638
rect -1006 -3774 -806 -3758
rect -1006 -3808 -990 -3774
rect -822 -3808 -806 -3774
rect -1006 -3831 -806 -3808
rect -1006 -4184 -806 -4161
rect -1006 -4218 -990 -4184
rect -822 -4218 -806 -4184
rect -1006 -4234 -806 -4218
<< polycont >>
rect -990 832 -822 866
rect -990 422 -822 456
rect -990 252 -822 286
rect -990 -158 -822 -124
rect -990 -328 -822 -294
rect -990 -738 -822 -704
rect -990 -908 -822 -874
rect -990 -1318 -822 -1284
rect -990 -1488 -822 -1454
rect -990 -1898 -822 -1864
rect -990 -2068 -822 -2034
rect -990 -2478 -822 -2444
rect -990 -2648 -822 -2614
rect -990 -3058 -822 -3024
rect -990 -3228 -822 -3194
rect -990 -3638 -822 -3604
rect -990 -3808 -822 -3774
rect -990 -4218 -822 -4184
<< npolyres >>
rect -1006 479 -806 809
rect -1006 -101 -806 229
rect -1006 -681 -806 -351
rect -1006 -1261 -806 -931
rect -1006 -1841 -806 -1511
rect -1006 -2421 -806 -2091
rect -1006 -3001 -806 -2671
rect -1006 -3581 -806 -3251
rect -1006 -4161 -806 -3831
<< locali >>
rect -1006 832 -990 866
rect -822 832 -806 866
rect -1006 422 -990 456
rect -822 422 -806 456
rect -1006 252 -990 286
rect -822 252 -806 286
rect -1006 -158 -990 -124
rect -822 -158 -806 -124
rect -1006 -328 -990 -294
rect -822 -328 -806 -294
rect -1006 -738 -990 -704
rect -822 -738 -806 -704
rect -1006 -908 -990 -874
rect -822 -908 -806 -874
rect -1006 -1318 -990 -1284
rect -822 -1318 -806 -1284
rect -1006 -1488 -990 -1454
rect -822 -1488 -806 -1454
rect -1006 -1898 -990 -1864
rect -822 -1898 -806 -1864
rect -1006 -2068 -990 -2034
rect -822 -2068 -806 -2034
rect -1006 -2478 -990 -2444
rect -822 -2478 -806 -2444
rect -1006 -2648 -990 -2614
rect -822 -2648 -806 -2614
rect -1006 -3058 -990 -3024
rect -822 -3058 -806 -3024
rect -1006 -3228 -990 -3194
rect -822 -3228 -806 -3194
rect -1006 -3638 -990 -3604
rect -822 -3638 -806 -3604
rect -1006 -3808 -990 -3774
rect -822 -3808 -806 -3774
rect -1006 -4218 -990 -4184
rect -822 -4218 -806 -4184
<< viali >>
rect -990 832 -822 866
rect -990 826 -822 832
rect -990 456 -822 462
rect -990 422 -822 456
rect -990 252 -822 286
rect -990 246 -822 252
rect -990 -124 -822 -118
rect -990 -158 -822 -124
rect -990 -328 -822 -294
rect -990 -334 -822 -328
rect -990 -704 -822 -698
rect -990 -738 -822 -704
rect -990 -908 -822 -874
rect -990 -914 -822 -908
rect -990 -1284 -822 -1278
rect -990 -1318 -822 -1284
rect -990 -1488 -822 -1454
rect -990 -1494 -822 -1488
rect -990 -1864 -822 -1858
rect -990 -1898 -822 -1864
rect -990 -2068 -822 -2034
rect -990 -2074 -822 -2068
rect -990 -2444 -822 -2438
rect -990 -2478 -822 -2444
rect -990 -2648 -822 -2614
rect -990 -2654 -822 -2648
rect -990 -3024 -822 -3018
rect -990 -3058 -822 -3024
rect -990 -3228 -822 -3194
rect -990 -3234 -822 -3228
rect -990 -3604 -822 -3598
rect -990 -3638 -822 -3604
rect -990 -3808 -822 -3774
rect -990 -3814 -822 -3808
rect -990 -4184 -822 -4178
rect -990 -4218 -822 -4184
<< metal1 >>
rect -1002 866 -810 872
rect -1002 826 -990 866
rect -822 826 -810 866
rect -1002 820 -810 826
rect -1002 462 -810 468
rect -1002 422 -990 462
rect -822 422 -810 462
rect -1002 416 -810 422
rect -1002 286 -810 292
rect -1002 246 -990 286
rect -822 246 -810 286
rect -1002 240 -810 246
rect -1002 -118 -810 -112
rect -1002 -158 -990 -118
rect -822 -158 -810 -118
rect -1002 -164 -810 -158
rect -1002 -294 -810 -288
rect -1002 -334 -990 -294
rect -822 -334 -810 -294
rect -1002 -340 -810 -334
rect -1002 -698 -810 -692
rect -1002 -738 -990 -698
rect -822 -738 -810 -698
rect -1002 -744 -810 -738
rect -1002 -874 -810 -868
rect -1002 -914 -990 -874
rect -822 -914 -810 -874
rect -1002 -920 -810 -914
rect -1002 -1278 -810 -1272
rect -1002 -1318 -990 -1278
rect -822 -1318 -810 -1278
rect -1002 -1324 -810 -1318
rect -1002 -1454 -810 -1448
rect -1002 -1494 -990 -1454
rect -822 -1494 -810 -1454
rect -1002 -1500 -810 -1494
rect -1002 -1858 -810 -1852
rect -1002 -1898 -990 -1858
rect -822 -1898 -810 -1858
rect -1002 -1904 -810 -1898
rect -1002 -2034 -810 -2028
rect -1002 -2074 -990 -2034
rect -822 -2074 -810 -2034
rect -1002 -2080 -810 -2074
rect -1002 -2438 -810 -2432
rect -1002 -2478 -990 -2438
rect -822 -2478 -810 -2438
rect -1002 -2484 -810 -2478
rect -1002 -2614 -810 -2608
rect -1002 -2654 -990 -2614
rect -822 -2654 -810 -2614
rect -1002 -2660 -810 -2654
rect -1002 -3018 -810 -3012
rect -1002 -3058 -990 -3018
rect -822 -3058 -810 -3018
rect -1002 -3064 -810 -3058
rect -1002 -3194 -810 -3188
rect -1002 -3234 -990 -3194
rect -822 -3234 -810 -3194
rect -1002 -3240 -810 -3234
rect -1002 -3598 -810 -3592
rect -1002 -3638 -990 -3598
rect -822 -3638 -810 -3598
rect -1002 -3644 -810 -3638
rect -1002 -3774 -810 -3768
rect -1002 -3814 -990 -3774
rect -822 -3814 -810 -3774
rect -1002 -3820 -810 -3814
rect -1002 -4178 -810 -4172
rect -1002 -4218 -990 -4178
rect -822 -4218 -810 -4178
rect -1002 -4224 -810 -4218
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 1 l 1.650 m 10 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 48.2 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 0 grc 0 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 0 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
