magic
tech sky130A
magscale 1 2
timestamp 1662126094
<< nwell >>
rect -209 -121 317 417
<< pmos >>
rect -9 98 21 198
rect 87 98 117 198
<< pdiff >>
rect -71 186 -9 198
rect -71 110 -59 186
rect -25 110 -9 186
rect -71 98 -9 110
rect 21 186 87 198
rect 21 110 37 186
rect 71 110 87 186
rect 21 98 87 110
rect 117 186 179 198
rect 117 110 133 186
rect 167 110 179 186
rect 117 98 179 110
<< pdiffc >>
rect -59 110 -25 186
rect 37 110 71 186
rect 133 110 167 186
<< nsubdiff >>
rect -173 347 -77 381
rect 185 347 281 381
rect -173 285 -139 347
rect 247 285 281 347
rect -173 -51 -139 11
rect 247 -51 281 11
rect -173 -85 -77 -51
rect 185 -85 281 -51
<< nsubdiffcont >>
rect -77 347 185 381
rect -173 11 -139 285
rect 247 11 281 285
rect -77 -85 185 -51
<< poly >>
rect 69 280 135 295
rect -9 279 135 280
rect -9 249 85 279
rect -9 198 21 249
rect 69 245 85 249
rect 119 245 135 279
rect 69 229 135 245
rect 87 198 117 229
rect -9 67 21 98
rect 87 72 117 98
<< polycont >>
rect 85 245 119 279
<< locali >>
rect -173 347 -77 381
rect 185 347 281 381
rect -173 285 -139 347
rect 247 285 281 347
rect 69 245 85 279
rect 119 245 135 279
rect -173 -51 -139 11
rect -59 186 -25 202
rect -59 44 -25 110
rect 37 186 71 202
rect 37 94 71 110
rect 133 186 167 202
rect 133 44 167 110
rect -59 10 167 44
rect -59 -51 -25 10
rect 247 -51 281 11
rect -173 -85 -77 -51
rect 185 -85 281 -51
rect -59 -553 -25 -85
rect -71 -573 -7 -553
rect -71 -608 -58 -573
rect -20 -608 -7 -573
rect -71 -625 -7 -608
<< viali >>
rect 85 245 119 279
rect -59 110 -25 186
rect 37 110 71 186
rect 133 110 167 186
rect -58 -608 -20 -573
<< metal1 >>
rect 3314 3986 7973 4089
rect 3314 3595 3417 3986
rect 3257 3363 3455 3595
rect 3256 2977 3454 3014
rect 3256 2858 7655 2977
rect 3256 2782 3454 2858
rect 3255 2378 3453 2435
rect 3255 2258 7419 2378
rect 3255 2203 3453 2258
rect 3256 1817 3454 1854
rect 3256 1687 7200 1817
rect 3256 1622 3454 1687
rect 7070 1285 7200 1687
rect 7299 1680 7419 2258
rect 7536 2080 7655 2858
rect 7870 2369 7973 3986
rect 7536 1961 7981 2080
rect 7299 1560 7981 1680
rect 3255 1217 3453 1273
rect 3255 1156 6754 1217
rect 1231 1122 6754 1156
rect 7070 1155 7986 1285
rect 73 279 131 285
rect 31 248 85 279
rect 69 245 85 248
rect 119 245 131 279
rect 1231 261 1265 1122
rect 3255 1085 6754 1122
rect 3255 1041 3453 1085
rect 6622 886 6754 1085
rect 6622 754 7987 886
rect 3255 653 3453 695
rect 3255 516 6226 653
rect 3255 463 3453 516
rect 6089 489 6226 516
rect 6089 352 7990 489
rect 73 239 131 245
rect 569 227 1274 261
rect -65 186 -19 198
rect -65 110 -59 186
rect -25 110 -19 186
rect -65 98 -19 110
rect 31 186 77 198
rect 31 110 37 186
rect 71 110 77 186
rect 31 98 77 110
rect 127 186 173 198
rect 127 110 133 186
rect 167 110 173 186
rect 127 98 173 110
rect 37 -251 71 98
rect 569 -251 603 227
rect 3258 89 3456 113
rect 3258 -48 7990 89
rect 3258 -119 3456 -48
rect 37 -285 603 -251
rect 4901 -458 7999 -302
rect 3257 -538 3455 -466
rect 4901 -538 5057 -458
rect -90 -573 -1 -547
rect -90 -608 -58 -573
rect -20 -608 -1 -573
rect -90 -627 -1 -608
rect -89 -906 -16 -627
rect 3257 -694 5057 -538
rect 3257 -698 3455 -694
rect 5235 -854 7995 -706
rect 3253 -1094 3451 -1037
rect 5235 -1094 5383 -854
rect 3253 -1242 5383 -1094
rect 3253 -1269 3451 -1242
rect 3255 -2209 3453 -1628
rect 5357 -1668 8003 -1533
rect 5357 -2209 5492 -1668
rect 3255 -2344 5492 -2209
<< properties >>
string FIXED_BBOX -210 -216 210 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
