magic
tech sky130A
magscale 1 2
timestamp 1662126094
<< poly >>
rect 3834 4172 4034 4188
rect 3834 4138 3850 4172
rect 4018 4138 4034 4172
rect 3834 4115 4034 4138
rect 3834 3762 4034 3785
rect 3834 3728 3850 3762
rect 4018 3728 4034 3762
rect 3834 3712 4034 3728
rect 3834 3592 4034 3608
rect 3834 3558 3850 3592
rect 4018 3558 4034 3592
rect 3834 3535 4034 3558
rect 3834 3182 4034 3205
rect 3834 3148 3850 3182
rect 4018 3148 4034 3182
rect 3834 3132 4034 3148
rect 3834 3012 4034 3028
rect 3834 2978 3850 3012
rect 4018 2978 4034 3012
rect 3834 2955 4034 2978
rect 3834 2602 4034 2625
rect 3834 2568 3850 2602
rect 4018 2568 4034 2602
rect 3834 2552 4034 2568
rect 3834 2432 4034 2448
rect 3834 2398 3850 2432
rect 4018 2398 4034 2432
rect 3834 2375 4034 2398
rect 3834 2022 4034 2045
rect 3834 1988 3850 2022
rect 4018 1988 4034 2022
rect 3834 1972 4034 1988
rect 3834 1852 4034 1868
rect 3834 1818 3850 1852
rect 4018 1818 4034 1852
rect 3834 1795 4034 1818
rect 3834 1442 4034 1465
rect 3834 1408 3850 1442
rect 4018 1408 4034 1442
rect 3834 1392 4034 1408
rect 3834 1272 4034 1288
rect 3834 1238 3850 1272
rect 4018 1238 4034 1272
rect 3834 1215 4034 1238
rect 3834 862 4034 885
rect 3834 828 3850 862
rect 4018 828 4034 862
rect 3834 812 4034 828
rect 3834 692 4034 708
rect 3834 658 3850 692
rect 4018 658 4034 692
rect 3834 635 4034 658
rect 3834 282 4034 305
rect 3834 248 3850 282
rect 4018 248 4034 282
rect 3834 232 4034 248
rect 3834 112 4034 128
rect 3834 78 3850 112
rect 4018 78 4034 112
rect 3834 55 4034 78
rect 3834 -298 4034 -275
rect 3834 -332 3850 -298
rect 4018 -332 4034 -298
rect 3834 -348 4034 -332
rect 3834 -468 4034 -452
rect 3834 -502 3850 -468
rect 4018 -502 4034 -468
rect 3834 -525 4034 -502
rect 3834 -878 4034 -855
rect 3834 -912 3850 -878
rect 4018 -912 4034 -878
rect 3834 -928 4034 -912
<< polycont >>
rect 3850 4138 4018 4172
rect 3850 3728 4018 3762
rect 3850 3558 4018 3592
rect 3850 3148 4018 3182
rect 3850 2978 4018 3012
rect 3850 2568 4018 2602
rect 3850 2398 4018 2432
rect 3850 1988 4018 2022
rect 3850 1818 4018 1852
rect 3850 1408 4018 1442
rect 3850 1238 4018 1272
rect 3850 828 4018 862
rect 3850 658 4018 692
rect 3850 248 4018 282
rect 3850 78 4018 112
rect 3850 -332 4018 -298
rect 3850 -502 4018 -468
rect 3850 -912 4018 -878
<< npolyres >>
rect 3834 3785 4034 4115
rect 3834 3205 4034 3535
rect 3834 2625 4034 2955
rect 3834 2045 4034 2375
rect 3834 1465 4034 1795
rect 3834 885 4034 1215
rect 3834 305 4034 635
rect 3834 -275 4034 55
rect 3834 -855 4034 -525
<< locali >>
rect 3834 4138 3850 4172
rect 4018 4138 4034 4172
rect 3834 3728 3850 3762
rect 4018 3728 4034 3762
rect 3834 3558 3850 3592
rect 4018 3558 4034 3592
rect 3834 3148 3850 3182
rect 4018 3148 4034 3182
rect 3834 2978 3850 3012
rect 4018 2978 4034 3012
rect 3834 2568 3850 2602
rect 4018 2568 4034 2602
rect 3834 2398 3850 2432
rect 4018 2398 4034 2432
rect 3834 1988 3850 2022
rect 4018 1988 4034 2022
rect 3834 1818 3850 1852
rect 4018 1818 4034 1852
rect 3834 1408 3850 1442
rect 4018 1408 4034 1442
rect 3834 1238 3850 1272
rect 4018 1238 4034 1272
rect 3834 828 3850 862
rect 4018 828 4034 862
rect 3834 658 3850 692
rect 4018 658 4034 692
rect 3834 248 3850 282
rect 4018 248 4034 282
rect 3834 78 3850 112
rect 4018 78 4034 112
rect 3834 -332 3850 -298
rect 4018 -332 4034 -298
rect 3834 -502 3850 -468
rect 4018 -502 4034 -468
rect 3834 -912 3850 -878
rect 4018 -912 4034 -878
<< viali >>
rect 3850 4138 4018 4172
rect 3850 4132 4018 4138
rect 3850 3762 4018 3768
rect 3850 3728 4018 3762
rect 3850 3558 4018 3592
rect 3850 3552 4018 3558
rect 3850 3182 4018 3188
rect 3850 3148 4018 3182
rect 3850 2978 4018 3012
rect 3850 2972 4018 2978
rect 3850 2602 4018 2608
rect 3850 2568 4018 2602
rect 3850 2398 4018 2432
rect 3850 2392 4018 2398
rect 3850 2022 4018 2028
rect 3850 1988 4018 2022
rect 3850 1818 4018 1852
rect 3850 1812 4018 1818
rect 3850 1442 4018 1448
rect 3850 1408 4018 1442
rect 3850 1238 4018 1272
rect 3850 1232 4018 1238
rect 3850 862 4018 868
rect 3850 828 4018 862
rect 3850 658 4018 692
rect 3850 652 4018 658
rect 3850 282 4018 288
rect 3850 248 4018 282
rect 3850 78 4018 112
rect 3850 72 4018 78
rect 3850 -298 4018 -292
rect 3850 -332 4018 -298
rect 3850 -502 4018 -468
rect 3850 -508 4018 -502
rect 3850 -878 4018 -872
rect 3850 -912 4018 -878
<< metal1 >>
rect 3838 4172 4030 4178
rect 3838 4132 3850 4172
rect 4018 4132 4030 4172
rect 3838 4126 4030 4132
rect 3838 3768 4030 3774
rect 3838 3728 3850 3768
rect 4018 3728 4030 3768
rect 3838 3722 4030 3728
rect 3838 3592 4030 3598
rect 3838 3552 3850 3592
rect 4018 3552 4030 3592
rect 3838 3546 4030 3552
rect -7667 3240 -7467 3440
rect 3838 3188 4030 3194
rect 3838 3148 3850 3188
rect 4018 3148 4030 3188
rect 3838 3142 4030 3148
rect 8400 3083 8600 3283
rect -7667 2840 -7467 3040
rect 3838 3012 4030 3018
rect 3838 2972 3850 3012
rect 4018 2972 4030 3012
rect 3838 2966 4030 2972
rect 8400 2683 8600 2883
rect -7667 2440 -7467 2640
rect 3838 2608 4030 2614
rect 3838 2568 3850 2608
rect 4018 2568 4030 2608
rect 3838 2562 4030 2568
rect 3838 2432 4030 2438
rect 3838 2392 3850 2432
rect 4018 2392 4030 2432
rect 3838 2386 4030 2392
rect 8400 2283 8600 2483
rect -7667 2040 -7467 2240
rect 3838 2028 4030 2034
rect 3838 1988 3850 2028
rect 4018 1988 4030 2028
rect 3838 1982 4030 1988
rect 8400 1883 8600 2083
rect 3838 1852 4030 1858
rect -7667 1640 -7467 1840
rect 3838 1812 3850 1852
rect 4018 1812 4030 1852
rect 3838 1806 4030 1812
rect 8400 1483 8600 1683
rect 3838 1448 4030 1454
rect -7667 1240 -7467 1440
rect 3838 1408 3850 1448
rect 4018 1408 4030 1448
rect 3838 1402 4030 1408
rect 3838 1272 4030 1278
rect 3838 1232 3850 1272
rect 4018 1232 4030 1272
rect 3838 1226 4030 1232
rect 8400 1083 8600 1283
rect -7667 840 -7467 1040
rect 3838 868 4030 874
rect 3838 828 3850 868
rect 4018 828 4030 868
rect 3838 822 4030 828
rect 3838 692 4030 698
rect 3838 652 3850 692
rect 4018 652 4030 692
rect 8400 683 8600 883
rect 3838 646 4030 652
rect -7667 440 -7467 640
rect 3838 288 4030 294
rect 3838 248 3850 288
rect 4018 248 4030 288
rect 8400 283 8600 483
rect 3838 242 4030 248
rect -7667 40 -7467 240
rect 3838 112 4030 118
rect 3838 72 3850 112
rect 4018 72 4030 112
rect 3838 66 4030 72
rect -7667 -360 -7467 -160
rect -664 -200 -464 0
rect 426 -207 626 -7
rect 8400 -117 8600 83
rect 3838 -292 4030 -286
rect 3838 -332 3850 -292
rect 4018 -332 4030 -292
rect 3838 -338 4030 -332
rect 3838 -468 4030 -462
rect 3838 -508 3850 -468
rect 4018 -508 4030 -468
rect 3838 -514 4030 -508
rect 3838 -872 4030 -866
rect 3838 -912 3850 -872
rect 4018 -912 4030 -872
rect 3838 -918 4030 -912
rect 8414 -938 8614 -738
use sky130_fd_pr__res_generic_po_4WEV9M  R1
timestamp 1662121956
transform 1 0 1055 0 1 845
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R2
timestamp 1662121956
transform 1 0 1534 0 1 792
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R3
timestamp 1662121956
transform 1 0 2013 0 1 739
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R4
timestamp 1662121956
transform 1 0 2492 0 1 686
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R5
timestamp 1662121956
transform 1 0 2971 0 1 633
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R6
timestamp 1662121956
transform 1 0 3450 0 1 580
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R7
timestamp 1662121956
transform 1 0 3929 0 1 527
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R8
timestamp 1662121956
transform 1 0 4408 0 1 474
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R9
timestamp 1662121956
transform 1 0 4887 0 1 421
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R10
timestamp 1662121956
transform 1 0 5366 0 1 368
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R11
timestamp 1662121956
transform 1 0 5845 0 1 315
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R12
timestamp 1662121956
transform 1 0 6324 0 1 262
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R13
timestamp 1662121956
transform 1 0 6803 0 1 209
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R14
timestamp 1662121956
transform 1 0 7282 0 1 156
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R15
timestamp 1662121956
transform 1 0 7761 0 1 103
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R16
timestamp 1662121956
transform 1 0 8240 0 1 50
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R17
timestamp 1662121956
transform 1 0 8719 0 1 -3
box 0 0 1 1
use sky130_fd_pr__res_generic_po_4WEV9M  R18
timestamp 1662121956
transform 1 0 9198 0 1 -56
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1662126094
transform 1 0 158 0 1 857
box -7819 -2633 631 3771
use sky130_fd_pr__pfet_01v8_XJT6XQ  XM2
timestamp 1662126094
transform 1 0 579 0 1 763
box -209 -2344 8003 4089
use sky130_fd_pr__res_generic_po_C4R5Y4  sky130_fd_pr__res_generic_po_C4R5Y4_0
timestamp 1662121956
transform 1 0 7201 0 1 2768
box 0 0 1 1
use sky130_fd_pr__res_generic_po_JD8CB6  sky130_fd_pr__res_generic_po_JD8CB6_0
timestamp 1662126094
transform 1 0 -2840 0 1 3010
box -1006 -4234 -806 882
<< labels >>
flabel metal1 -664 -200 -464 0 0 FreeSans 256 0 0 0 VN
port 10 nsew
flabel metal1 426 -207 626 -7 0 FreeSans 256 0 0 0 VP
port 9 nsew
flabel metal1 8400 3083 8600 3283 0 FreeSans 256 0 0 0 Y0
port 0 nsew
flabel metal1 8400 2683 8600 2883 0 FreeSans 256 0 0 0 Y1
port 1 nsew
flabel metal1 8400 2283 8600 2483 0 FreeSans 256 0 0 0 Y2
port 2 nsew
flabel metal1 8400 1883 8600 2083 0 FreeSans 256 0 0 0 Y3
port 3 nsew
flabel metal1 8400 1483 8600 1683 0 FreeSans 256 0 0 0 Y4
port 4 nsew
flabel metal1 8400 1083 8600 1283 0 FreeSans 256 0 0 0 Y5
port 5 nsew
flabel metal1 8400 683 8600 883 0 FreeSans 256 0 0 0 Y6
port 6 nsew
flabel metal1 8400 283 8600 483 0 FreeSans 256 0 0 0 Y7
port 7 nsew
flabel metal1 8400 -117 8600 83 0 FreeSans 256 0 0 0 Y8
port 8 nsew
flabel metal1 8414 -938 8614 -738 0 FreeSans 256 0 0 0 Y9
port 21 nsew
flabel metal1 -7667 3240 -7467 3440 0 FreeSans 256 0 0 0 I0
port 20 nsew
flabel metal1 -7667 2840 -7467 3040 0 FreeSans 256 0 0 0 I1
port 19 nsew
flabel metal1 -7667 2440 -7467 2640 0 FreeSans 256 0 0 0 I2
port 18 nsew
flabel metal1 -7667 2040 -7467 2240 0 FreeSans 256 0 0 0 I3
port 17 nsew
flabel metal1 -7667 1640 -7467 1840 0 FreeSans 256 0 0 0 I4
port 16 nsew
flabel metal1 -7667 1240 -7467 1440 0 FreeSans 256 0 0 0 I5
port 15 nsew
flabel metal1 -7667 840 -7467 1040 0 FreeSans 256 0 0 0 I6
port 14 nsew
flabel metal1 -7667 440 -7467 640 0 FreeSans 256 0 0 0 I7
port 13 nsew
flabel metal1 -7667 40 -7467 240 0 FreeSans 256 0 0 0 I8
port 12 nsew
flabel metal1 -7667 -360 -7467 -160 0 FreeSans 256 0 0 0 I9
port 11 nsew
<< end >>
